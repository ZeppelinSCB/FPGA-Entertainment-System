module letter_snake_game
(
    letter_x        ,
    letter_y        ,
    letter_press    ,
    letter_press_o        
);

input   [7:0]   letter_x     ;//x coordinate of pixel with respect to letter
input   [7:0]   letter_y     ;//y coordinate of pixel with respect to letter

output  [0:0]   letter_o     ;//letter output


assign          letter_press[ 0] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_press[ 1] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_press[ 2] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_press[ 3] <= {8'b11111100, 8'b00000000, 8'b11111100, 8'b00000000, 8'b11111100, 8'b00000000, 8'b00111110, 8'b00000000, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00010000, 8'b00000000, 8'b11000111, 8'b00000000, 8'b11101110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11101110, 8'b00000000, 8'b11111100, 8'b00000000, 8'b11101110, 8'b00000000};
assign          letter_press[ 4] <= {8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00010000, 8'b00000000, 8'b01100010, 8'b00000000, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000100, 8'b00000000};
assign          letter_press[ 5] <= {8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01001000, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011000, 8'b00000000, 8'b01100010, 8'b00000000, 8'b01000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b01000100, 8'b00000000};
assign          letter_press[ 6] <= {8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01001000, 8'b00000000, 8'b01000000, 8'b00000000, 8'b01000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101000, 8'b00000000, 8'b01010010, 8'b00000000, 8'b00101000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01010000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b00101000, 8'b00000000};
assign          letter_press[ 7] <= {8'b01000010, 8'b00000000, 8'b01111100, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00100000, 8'b00000000, 8'b00100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00101000, 8'b00000000, 8'b01010010, 8'b00000000, 8'b00101000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00101000, 8'b00000000};
assign          letter_press[ 8] <= {8'b01111100, 8'b00000000, 8'b01001000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b00011000, 8'b00000000, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00100100, 8'b00000000, 8'b01001010, 8'b00000000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01010000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b00010000, 8'b00000000};
assign          letter_press[ 9] <= {8'b01000000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000000, 8'b01001010, 8'b00000000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b00010000, 8'b00000000};
assign          letter_press[10] <= {8'b01000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b01000000, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b01001010, 8'b00000000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01001000, 8'b00000000, 8'b01000000, 8'b00000000, 8'b00010000, 8'b00000000};
assign          letter_press[11] <= {8'b01000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000110, 8'b00000000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b01000010, 8'b00000000, 8'b00010000, 8'b00000000};
assign          letter_press[12] <= {8'b01000000, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000010, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000010, 8'b00000000, 8'b01000110, 8'b00000000, 8'b00010000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01000100, 8'b00000000, 8'b01000010, 8'b00000000, 8'b00010000, 8'b00000000};
assign          letter_press[13] <= {8'b11100000, 8'b00000000, 8'b11100011, 8'b00000000, 8'b11111100, 8'b00000000, 8'b01111100, 8'b00000000, 8'b01111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11100111, 8'b00000000, 8'b11100010, 8'b00000000, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11101110, 8'b00000000, 8'b11111100, 8'b00000000, 8'b00111000, 8'b00000000};
assign          letter_press[14] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_press[15] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};

always@(*)
begin
    letter_press_o = letter[letter_y][letter_x];
end

endmodule