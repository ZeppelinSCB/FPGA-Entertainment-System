module letter_game_over
(
    letter_x        ,
    letter_y        ,
    letter_over    ,
    letter_over_o        
);

input   [7:0]   letter_x     ;//x coordinate of pixel with respect to letter
input   [7:0]   letter_y     ;//y coordinate of pixel with respect to letter

output  [0:0]   letter_over_o     ;//letter output


assign          letter_over[ 0] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[ 1] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[ 2] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[ 3] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[ 4] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[ 5] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[ 6] <= {8'b00000000, 8'b11111110, 8'b01111111, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11100000, 8'b00000000};
assign          letter_over[ 7] <= {8'b00000000, 8'b01111100, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b01111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111101, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01111110, 8'b00000000, 8'b00000000, 8'b01111101, 8'b11111000, 8'b00000000};
assign          letter_over[ 8] <= {8'b00000000, 8'b00111100, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b01111100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b01111100, 8'b00000000};
assign          letter_over[ 9] <= {8'b00000000, 8'b00111100, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011100, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00111100, 8'b00000000};
assign          letter_over[10] <= {8'b00000000, 8'b00011100, 8'b00111000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_over[11] <= {8'b00000000, 8'b00011110, 8'b00111000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_over[12] <= {8'b00000000, 8'b00011110, 8'b01110000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_over[13] <= {8'b00000000, 8'b00001111, 8'b01110000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001110, 8'b00000000};
assign          letter_over[14] <= {8'b00000000, 8'b00001111, 8'b01100000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_over[15] <= {8'b00000000, 8'b00001111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_over[16] <= {8'b00000000, 8'b00000111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_over[17] <= {8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_over[18] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_over[19] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_over[20] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_over[21] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_over[22] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000011, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_over[23] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_over[24] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00111100, 8'b00000000};
assign          letter_over[25] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b01111000, 8'b00000000};
assign          letter_over[26] <= {8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01111110, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11111000, 8'b00000000};
assign          letter_over[27] <= {8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11100000, 8'b00000000};
assign          letter_over[28] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[29] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[30] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_over[31] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};


always@(*)
begin
    letter_over_o = letter_over[letter_y][letter_x];
end

endmodule