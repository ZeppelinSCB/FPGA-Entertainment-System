`include "../libs/define.vh"

module start_page
(
    vga_clk,
    sys_rst_n,
    clk
);



endmodule