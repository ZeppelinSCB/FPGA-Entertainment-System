`include "../libs/define.vh"

module start_page
(
    vga_clk,
    sys_rst_n,
    one_resistor_x,
    two_resistors_x,
    one_resistor_y,
    two_resistors_y,
    clk
);



endmodule