`ifndef sprites_vh
`define sprites_vh

`define APPLE_PIC \
sp[4'd8][0][0] = 3'b111;\
sp[4'd8][0][1] = 3'b111;\
sp[4'd8][0][2] = 3'b111;\
sp[4'd8][0][3] = 3'b111;\
sp[4'd8][0][4] = 3'b111;\
sp[4'd8][0][5] = 3'b111;\
sp[4'd8][0][6] = 3'b111;\
sp[4'd8][0][7] = 3'b111;\
sp[4'd8][0][8] = 3'b111;\
sp[4'd8][0][9] = 3'b111;\
sp[4'd8][0][10] = 3'b111;\
sp[4'd8][0][11] = 3'b111;\
sp[4'd8][0][12] = 3'b111;\
sp[4'd8][0][13] = 3'b111;\
sp[4'd8][0][14] = 3'b111;\
sp[4'd8][0][15] = 3'b111;\
sp[4'd8][1][0] = 3'b111;\
sp[4'd8][1][1] = 3'b111;\
sp[4'd8][1][2] = 3'b111;\
sp[4'd8][1][3] = 3'b111;\
sp[4'd8][1][4] = 3'b111;\
sp[4'd8][1][5] = 3'b111;\
sp[4'd8][1][6] = 3'b111;\
sp[4'd8][1][7] = 3'b111;\
sp[4'd8][1][8] = 3'b111;\
sp[4'd8][1][9] = 3'b111;\
sp[4'd8][1][10] = 3'b111;\
sp[4'd8][1][11] = 3'b111;\
sp[4'd8][1][12] = 3'b111;\
sp[4'd8][1][13] = 3'b111;\
sp[4'd8][1][14] = 3'b111;\
sp[4'd8][1][15] = 3'b111;\
sp[4'd8][2][0] = 3'b111;\
sp[4'd8][2][1] = 3'b111;\
sp[4'd8][2][2] = 3'b111;\
sp[4'd8][2][3] = 3'b111;\
sp[4'd8][2][4] = 3'b111;\
sp[4'd8][2][5] = 3'b111;\
sp[4'd8][2][6] = 3'b111;\
sp[4'd8][2][7] = 3'b111;\
sp[4'd8][2][8] = 3'b111;\
sp[4'd8][2][9] = 3'b111;\
sp[4'd8][2][10] = 3'b111;\
sp[4'd8][2][11] = 3'b111;\
sp[4'd8][2][12] = 3'b111;\
sp[4'd8][2][13] = 3'b111;\
sp[4'd8][2][14] = 3'b111;\
sp[4'd8][2][15] = 3'b111;\
sp[4'd8][3][0] = 3'b111;\
sp[4'd8][3][1] = 3'b111;\
sp[4'd8][3][2] = 3'b111;\
sp[4'd8][3][3] = 3'b111;\
sp[4'd8][3][4] = 3'b111;\
sp[4'd8][3][5] = 3'b000;\
sp[4'd8][3][6] = 3'b000;\
sp[4'd8][3][7] = 3'b000;\
sp[4'd8][3][8] = 3'b000;\
sp[4'd8][3][9] = 3'b000;\
sp[4'd8][3][10] = 3'b000;\
sp[4'd8][3][11] = 3'b000;\
sp[4'd8][3][12] = 3'b000;\
sp[4'd8][3][13] = 3'b000;\
sp[4'd8][3][14] = 3'b111;\
sp[4'd8][3][15] = 3'b111;\
sp[4'd8][4][0] = 3'b111;\
sp[4'd8][4][1] = 3'b111;\
sp[4'd8][4][2] = 3'b111;\
sp[4'd8][4][3] = 3'b111;\
sp[4'd8][4][4] = 3'b000;\
sp[4'd8][4][5] = 3'b000;\
sp[4'd8][4][6] = 3'b100;\
sp[4'd8][4][7] = 3'b100;\
sp[4'd8][4][8] = 3'b100;\
sp[4'd8][4][9] = 3'b100;\
sp[4'd8][4][10] = 3'b100;\
sp[4'd8][4][11] = 3'b100;\
sp[4'd8][4][12] = 3'b100;\
sp[4'd8][4][13] = 3'b000;\
sp[4'd8][4][14] = 3'b000;\
sp[4'd8][4][15] = 3'b111;\
sp[4'd8][5][0] = 3'b111;\
sp[4'd8][5][1] = 3'b111;\
sp[4'd8][5][2] = 3'b111;\
sp[4'd8][5][3] = 3'b111;\
sp[4'd8][5][4] = 3'b000;\
sp[4'd8][5][5] = 3'b100;\
sp[4'd8][5][6] = 3'b100;\
sp[4'd8][5][7] = 3'b111;\
sp[4'd8][5][8] = 3'b111;\
sp[4'd8][5][9] = 3'b100;\
sp[4'd8][5][10] = 3'b100;\
sp[4'd8][5][11] = 3'b100;\
sp[4'd8][5][12] = 3'b100;\
sp[4'd8][5][13] = 3'b100;\
sp[4'd8][5][14] = 3'b000;\
sp[4'd8][5][15] = 3'b111;\
sp[4'd8][6][0] = 3'b111;\
sp[4'd8][6][1] = 3'b111;\
sp[4'd8][6][2] = 3'b111;\
sp[4'd8][6][3] = 3'b111;\
sp[4'd8][6][4] = 3'b000;\
sp[4'd8][6][5] = 3'b100;\
sp[4'd8][6][6] = 3'b100;\
sp[4'd8][6][7] = 3'b100;\
sp[4'd8][6][8] = 3'b100;\
sp[4'd8][6][9] = 3'b100;\
sp[4'd8][6][10] = 3'b100;\
sp[4'd8][6][11] = 3'b100;\
sp[4'd8][6][12] = 3'b100;\
sp[4'd8][6][13] = 3'b100;\
sp[4'd8][6][14] = 3'b000;\
sp[4'd8][6][15] = 3'b111;\
sp[4'd8][7][0] = 3'b111;\
sp[4'd8][7][1] = 3'b111;\
sp[4'd8][7][2] = 3'b111;\
sp[4'd8][7][3] = 3'b111;\
sp[4'd8][7][4] = 3'b000;\
sp[4'd8][7][5] = 3'b100;\
sp[4'd8][7][6] = 3'b000;\
sp[4'd8][7][7] = 3'b100;\
sp[4'd8][7][8] = 3'b100;\
sp[4'd8][7][9] = 3'b100;\
sp[4'd8][7][10] = 3'b100;\
sp[4'd8][7][11] = 3'b100;\
sp[4'd8][7][12] = 3'b100;\
sp[4'd8][7][13] = 3'b100;\
sp[4'd8][7][14] = 3'b000;\
sp[4'd8][7][15] = 3'b111;\
sp[4'd8][8][0] = 3'b111;\
sp[4'd8][8][1] = 3'b111;\
sp[4'd8][8][2] = 3'b000;\
sp[4'd8][8][3] = 3'b000;\
sp[4'd8][8][4] = 3'b000;\
sp[4'd8][8][5] = 3'b000;\
sp[4'd8][8][6] = 3'b000;\
sp[4'd8][8][7] = 3'b100;\
sp[4'd8][8][8] = 3'b100;\
sp[4'd8][8][9] = 3'b100;\
sp[4'd8][8][10] = 3'b100;\
sp[4'd8][8][11] = 3'b100;\
sp[4'd8][8][12] = 3'b100;\
sp[4'd8][8][13] = 3'b100;\
sp[4'd8][8][14] = 3'b000;\
sp[4'd8][8][15] = 3'b111;\
sp[4'd8][9][0] = 3'b111;\
sp[4'd8][9][1] = 3'b000;\
sp[4'd8][9][2] = 3'b000;\
sp[4'd8][9][3] = 3'b010;\
sp[4'd8][9][4] = 3'b010;\
sp[4'd8][9][5] = 3'b100;\
sp[4'd8][9][6] = 3'b000;\
sp[4'd8][9][7] = 3'b100;\
sp[4'd8][9][8] = 3'b100;\
sp[4'd8][9][9] = 3'b100;\
sp[4'd8][9][10] = 3'b100;\
sp[4'd8][9][11] = 3'b100;\
sp[4'd8][9][12] = 3'b100;\
sp[4'd8][9][13] = 3'b100;\
sp[4'd8][9][14] = 3'b000;\
sp[4'd8][9][15] = 3'b111;\
sp[4'd8][10][0] = 3'b111;\
sp[4'd8][10][1] = 3'b000;\
sp[4'd8][10][2] = 3'b010;\
sp[4'd8][10][3] = 3'b010;\
sp[4'd8][10][4] = 3'b010;\
sp[4'd8][10][5] = 3'b100;\
sp[4'd8][10][6] = 3'b100;\
sp[4'd8][10][7] = 3'b100;\
sp[4'd8][10][8] = 3'b100;\
sp[4'd8][10][9] = 3'b100;\
sp[4'd8][10][10] = 3'b100;\
sp[4'd8][10][11] = 3'b100;\
sp[4'd8][10][12] = 3'b100;\
sp[4'd8][10][13] = 3'b100;\
sp[4'd8][10][14] = 3'b000;\
sp[4'd8][10][15] = 3'b111;\
sp[4'd8][11][0] = 3'b111;\
sp[4'd8][11][1] = 3'b000;\
sp[4'd8][11][2] = 3'b010;\
sp[4'd8][11][3] = 3'b010;\
sp[4'd8][11][4] = 3'b000;\
sp[4'd8][11][5] = 3'b100;\
sp[4'd8][11][6] = 3'b100;\
sp[4'd8][11][7] = 3'b100;\
sp[4'd8][11][8] = 3'b100;\
sp[4'd8][11][9] = 3'b100;\
sp[4'd8][11][10] = 3'b100;\
sp[4'd8][11][11] = 3'b100;\
sp[4'd8][11][12] = 3'b100;\
sp[4'd8][11][13] = 3'b100;\
sp[4'd8][11][14] = 3'b000;\
sp[4'd8][11][15] = 3'b111;\
sp[4'd8][12][0] = 3'b111;\
sp[4'd8][12][1] = 3'b000;\
sp[4'd8][12][2] = 3'b000;\
sp[4'd8][12][3] = 3'b000;\
sp[4'd8][12][4] = 3'b000;\
sp[4'd8][12][5] = 3'b000;\
sp[4'd8][12][6] = 3'b100;\
sp[4'd8][12][7] = 3'b100;\
sp[4'd8][12][8] = 3'b100;\
sp[4'd8][12][9] = 3'b100;\
sp[4'd8][12][10] = 3'b100;\
sp[4'd8][12][11] = 3'b100;\
sp[4'd8][12][12] = 3'b100;\
sp[4'd8][12][13] = 3'b000;\
sp[4'd8][12][14] = 3'b000;\
sp[4'd8][12][15] = 3'b111;\
sp[4'd8][13][0] = 3'b111;\
sp[4'd8][13][1] = 3'b111;\
sp[4'd8][13][2] = 3'b111;\
sp[4'd8][13][3] = 3'b111;\
sp[4'd8][13][4] = 3'b111;\
sp[4'd8][13][5] = 3'b000;\
sp[4'd8][13][6] = 3'b000;\
sp[4'd8][13][7] = 3'b000;\
sp[4'd8][13][8] = 3'b000;\
sp[4'd8][13][9] = 3'b000;\
sp[4'd8][13][10] = 3'b000;\
sp[4'd8][13][11] = 3'b000;\
sp[4'd8][13][12] = 3'b000;\
sp[4'd8][13][13] = 3'b000;\
sp[4'd8][13][14] = 3'b111;\
sp[4'd8][13][15] = 3'b111;\
sp[4'd8][14][0] = 3'b111;\
sp[4'd8][14][1] = 3'b111;\
sp[4'd8][14][2] = 3'b111;\
sp[4'd8][14][3] = 3'b111;\
sp[4'd8][14][4] = 3'b111;\
sp[4'd8][14][5] = 3'b111;\
sp[4'd8][14][6] = 3'b111;\
sp[4'd8][14][7] = 3'b111;\
sp[4'd8][14][8] = 3'b111;\
sp[4'd8][14][9] = 3'b111;\
sp[4'd8][14][10] = 3'b111;\
sp[4'd8][14][11] = 3'b111;\
sp[4'd8][14][12] = 3'b111;\
sp[4'd8][14][13] = 3'b111;\
sp[4'd8][14][14] = 3'b111;\
sp[4'd8][14][15] = 3'b111;\
sp[4'd8][15][0] = 3'b111;\
sp[4'd8][15][1] = 3'b111;\
sp[4'd8][15][2] = 3'b111;\
sp[4'd8][15][3] = 3'b111;\
sp[4'd8][15][4] = 3'b111;\
sp[4'd8][15][5] = 3'b111;\
sp[4'd8][15][6] = 3'b111;\
sp[4'd8][15][7] = 3'b111;\
sp[4'd8][15][8] = 3'b111;\
sp[4'd8][15][9] = 3'b111;\
sp[4'd8][15][10] = 3'b111;\
sp[4'd8][15][11] = 3'b111;\
sp[4'd8][15][12] = 3'b111;\
sp[4'd8][15][13] = 3'b111;\
sp[4'd8][15][14] = 3'b111;\
sp[4'd8][15][15] = 3'b111;

`define SNAKE_HEAD_PIC \
sp[4'd4][0][0] = 3'b111;\
sp[4'd4][0][1] = 3'b111;\
sp[4'd4][0][2] = 3'b111;\
sp[4'd4][0][3] = 3'b111;\
sp[4'd4][0][4] = 3'b111;\
sp[4'd4][0][5] = 3'b111;\
sp[4'd4][0][6] = 3'b111;\
sp[4'd4][0][7] = 3'b111;\
sp[4'd4][0][8] = 3'b111;\
sp[4'd4][0][9] = 3'b111;\
sp[4'd4][0][10] = 3'b111;\
sp[4'd4][0][11] = 3'b111;\
sp[4'd4][0][12] = 3'b111;\
sp[4'd4][0][13] = 3'b111;\
sp[4'd4][0][14] = 3'b111;\
sp[4'd4][0][15] = 3'b111;\
sp[4'd4][1][0] = 3'b111;\
sp[4'd4][1][1] = 3'b111;\
sp[4'd4][1][2] = 3'b111;\
sp[4'd4][1][3] = 3'b111;\
sp[4'd4][1][4] = 3'b000;\
sp[4'd4][1][5] = 3'b000;\
sp[4'd4][1][6] = 3'b000;\
sp[4'd4][1][7] = 3'b000;\
sp[4'd4][1][8] = 3'b000;\
sp[4'd4][1][9] = 3'b000;\
sp[4'd4][1][10] = 3'b000;\
sp[4'd4][1][11] = 3'b111;\
sp[4'd4][1][12] = 3'b111;\
sp[4'd4][1][13] = 3'b111;\
sp[4'd4][1][14] = 3'b111;\
sp[4'd4][1][15] = 3'b111;\
sp[4'd4][2][0] = 3'b111;\
sp[4'd4][2][1] = 3'b111;\
sp[4'd4][2][2] = 3'b000;\
sp[4'd4][2][3] = 3'b000;\
sp[4'd4][2][4] = 3'b000;\
sp[4'd4][2][5] = 3'b010;\
sp[4'd4][2][6] = 3'b010;\
sp[4'd4][2][7] = 3'b010;\
sp[4'd4][2][8] = 3'b010;\
sp[4'd4][2][9] = 3'b010;\
sp[4'd4][2][10] = 3'b000;\
sp[4'd4][2][11] = 3'b000;\
sp[4'd4][2][12] = 3'b000;\
sp[4'd4][2][13] = 3'b111;\
sp[4'd4][2][14] = 3'b111;\
sp[4'd4][2][15] = 3'b111;\
sp[4'd4][3][0] = 3'b111;\
sp[4'd4][3][1] = 3'b000;\
sp[4'd4][3][2] = 3'b010;\
sp[4'd4][3][3] = 3'b010;\
sp[4'd4][3][4] = 3'b010;\
sp[4'd4][3][5] = 3'b010;\
sp[4'd4][3][6] = 3'b010;\
sp[4'd4][3][7] = 3'b010;\
sp[4'd4][3][8] = 3'b110;\
sp[4'd4][3][9] = 3'b010;\
sp[4'd4][3][10] = 3'b010;\
sp[4'd4][3][11] = 3'b010;\
sp[4'd4][3][12] = 3'b000;\
sp[4'd4][3][13] = 3'b000;\
sp[4'd4][3][14] = 3'b000;\
sp[4'd4][3][15] = 3'b111;\
sp[4'd4][4][0] = 3'b000;\
sp[4'd4][4][1] = 3'b010;\
sp[4'd4][4][2] = 3'b010;\
sp[4'd4][4][3] = 3'b111;\
sp[4'd4][4][4] = 3'b111;\
sp[4'd4][4][5] = 3'b111;\
sp[4'd4][4][6] = 3'b111;\
sp[4'd4][4][7] = 3'b010;\
sp[4'd4][4][8] = 3'b010;\
sp[4'd4][4][9] = 3'b010;\
sp[4'd4][4][10] = 3'b110;\
sp[4'd4][4][11] = 3'b010;\
sp[4'd4][4][12] = 3'b010;\
sp[4'd4][4][13] = 3'b010;\
sp[4'd4][4][14] = 3'b000;\
sp[4'd4][4][15] = 3'b000;\
sp[4'd4][5][0] = 3'b000;\
sp[4'd4][5][1] = 3'b010;\
sp[4'd4][5][2] = 3'b110;\
sp[4'd4][5][3] = 3'b111;\
sp[4'd4][5][4] = 3'b000;\
sp[4'd4][5][5] = 3'b000;\
sp[4'd4][5][6] = 3'b111;\
sp[4'd4][5][7] = 3'b010;\
sp[4'd4][5][8] = 3'b010;\
sp[4'd4][5][9] = 3'b010;\
sp[4'd4][5][10] = 3'b010;\
sp[4'd4][5][11] = 3'b010;\
sp[4'd4][5][12] = 3'b010;\
sp[4'd4][5][13] = 3'b110;\
sp[4'd4][5][14] = 3'b010;\
sp[4'd4][5][15] = 3'b000;\
sp[4'd4][6][0] = 3'b000;\
sp[4'd4][6][1] = 3'b110;\
sp[4'd4][6][2] = 3'b110;\
sp[4'd4][6][3] = 3'b111;\
sp[4'd4][6][4] = 3'b111;\
sp[4'd4][6][5] = 3'b111;\
sp[4'd4][6][6] = 3'b111;\
sp[4'd4][6][7] = 3'b010;\
sp[4'd4][6][8] = 3'b110;\
sp[4'd4][6][9] = 3'b010;\
sp[4'd4][6][10] = 3'b100;\
sp[4'd4][6][11] = 3'b010;\
sp[4'd4][6][12] = 3'b010;\
sp[4'd4][6][13] = 3'b010;\
sp[4'd4][6][14] = 3'b010;\
sp[4'd4][6][15] = 3'b000;\
sp[4'd4][7][0] = 3'b000;\
sp[4'd4][7][1] = 3'b010;\
sp[4'd4][7][2] = 3'b110;\
sp[4'd4][7][3] = 3'b010;\
sp[4'd4][7][4] = 3'b010;\
sp[4'd4][7][5] = 3'b010;\
sp[4'd4][7][6] = 3'b010;\
sp[4'd4][7][7] = 3'b010;\
sp[4'd4][7][8] = 3'b010;\
sp[4'd4][7][9] = 3'b010;\
sp[4'd4][7][10] = 3'b100;\
sp[4'd4][7][11] = 3'b010;\
sp[4'd4][7][12] = 3'b100;\
sp[4'd4][7][13] = 3'b010;\
sp[4'd4][7][14] = 3'b100;\
sp[4'd4][7][15] = 3'b000;\
sp[4'd4][8][0] = 3'b000;\
sp[4'd4][8][1] = 3'b010;\
sp[4'd4][8][2] = 3'b110;\
sp[4'd4][8][3] = 3'b010;\
sp[4'd4][8][4] = 3'b010;\
sp[4'd4][8][5] = 3'b010;\
sp[4'd4][8][6] = 3'b010;\
sp[4'd4][8][7] = 3'b110;\
sp[4'd4][8][8] = 3'b010;\
sp[4'd4][8][9] = 3'b010;\
sp[4'd4][8][10] = 3'b100;\
sp[4'd4][8][11] = 3'b100;\
sp[4'd4][8][12] = 3'b010;\
sp[4'd4][8][13] = 3'b100;\
sp[4'd4][8][14] = 3'b010;\
sp[4'd4][8][15] = 3'b000;\
sp[4'd4][9][0] = 3'b000;\
sp[4'd4][9][1] = 3'b110;\
sp[4'd4][9][2] = 3'b110;\
sp[4'd4][9][3] = 3'b111;\
sp[4'd4][9][4] = 3'b111;\
sp[4'd4][9][5] = 3'b111;\
sp[4'd4][9][6] = 3'b111;\
sp[4'd4][9][7] = 3'b010;\
sp[4'd4][9][8] = 3'b010;\
sp[4'd4][9][9] = 3'b010;\
sp[4'd4][9][10] = 3'b100;\
sp[4'd4][9][11] = 3'b010;\
sp[4'd4][9][12] = 3'b010;\
sp[4'd4][9][13] = 3'b010;\
sp[4'd4][9][14] = 3'b010;\
sp[4'd4][9][15] = 3'b000;\
sp[4'd4][10][0] = 3'b000;\
sp[4'd4][10][1] = 3'b010;\
sp[4'd4][10][2] = 3'b110;\
sp[4'd4][10][3] = 3'b111;\
sp[4'd4][10][4] = 3'b000;\
sp[4'd4][10][5] = 3'b000;\
sp[4'd4][10][6] = 3'b111;\
sp[4'd4][10][7] = 3'b010;\
sp[4'd4][10][8] = 3'b110;\
sp[4'd4][10][9] = 3'b010;\
sp[4'd4][10][10] = 3'b010;\
sp[4'd4][10][11] = 3'b010;\
sp[4'd4][10][12] = 3'b010;\
sp[4'd4][10][13] = 3'b010;\
sp[4'd4][10][14] = 3'b010;\
sp[4'd4][10][15] = 3'b000;\
sp[4'd4][11][0] = 3'b000;\
sp[4'd4][11][1] = 3'b010;\
sp[4'd4][11][2] = 3'b010;\
sp[4'd4][11][3] = 3'b111;\
sp[4'd4][11][4] = 3'b111;\
sp[4'd4][11][5] = 3'b111;\
sp[4'd4][11][6] = 3'b111;\
sp[4'd4][11][7] = 3'b010;\
sp[4'd4][11][8] = 3'b010;\
sp[4'd4][11][9] = 3'b010;\
sp[4'd4][11][10] = 3'b110;\
sp[4'd4][11][11] = 3'b010;\
sp[4'd4][11][12] = 3'b110;\
sp[4'd4][11][13] = 3'b010;\
sp[4'd4][11][14] = 3'b000;\
sp[4'd4][11][15] = 3'b000;\
sp[4'd4][12][0] = 3'b111;\
sp[4'd4][12][1] = 3'b000;\
sp[4'd4][12][2] = 3'b010;\
sp[4'd4][12][3] = 3'b010;\
sp[4'd4][12][4] = 3'b010;\
sp[4'd4][12][5] = 3'b010;\
sp[4'd4][12][6] = 3'b010;\
sp[4'd4][12][7] = 3'b010;\
sp[4'd4][12][8] = 3'b110;\
sp[4'd4][12][9] = 3'b010;\
sp[4'd4][12][10] = 3'b010;\
sp[4'd4][12][11] = 3'b010;\
sp[4'd4][12][12] = 3'b000;\
sp[4'd4][12][13] = 3'b000;\
sp[4'd4][12][14] = 3'b111;\
sp[4'd4][12][15] = 3'b111;\
sp[4'd4][13][0] = 3'b111;\
sp[4'd4][13][1] = 3'b111;\
sp[4'd4][13][2] = 3'b000;\
sp[4'd4][13][3] = 3'b000;\
sp[4'd4][13][4] = 3'b000;\
sp[4'd4][13][5] = 3'b010;\
sp[4'd4][13][6] = 3'b010;\
sp[4'd4][13][7] = 3'b010;\
sp[4'd4][13][8] = 3'b010;\
sp[4'd4][13][9] = 3'b010;\
sp[4'd4][13][10] = 3'b000;\
sp[4'd4][13][11] = 3'b000;\
sp[4'd4][13][12] = 3'b000;\
sp[4'd4][13][13] = 3'b111;\
sp[4'd4][13][14] = 3'b111;\
sp[4'd4][13][15] = 3'b111;\
sp[4'd4][14][0] = 3'b111;\
sp[4'd4][14][1] = 3'b111;\
sp[4'd4][14][2] = 3'b111;\
sp[4'd4][14][3] = 3'b111;\
sp[4'd4][14][4] = 3'b111;\
sp[4'd4][14][5] = 3'b000;\
sp[4'd4][14][6] = 3'b000;\
sp[4'd4][14][7] = 3'b000;\
sp[4'd4][14][8] = 3'b000;\
sp[4'd4][14][9] = 3'b000;\
sp[4'd4][14][10] = 3'b000;\
sp[4'd4][14][11] = 3'b111;\
sp[4'd4][14][12] = 3'b111;\
sp[4'd4][14][13] = 3'b111;\
sp[4'd4][14][14] = 3'b111;\
sp[4'd4][14][15] = 3'b111;\
sp[4'd4][15][0] = 3'b111;\
sp[4'd4][15][1] = 3'b111;\
sp[4'd4][15][2] = 3'b111;\
sp[4'd4][15][3] = 3'b111;\
sp[4'd4][15][4] = 3'b111;\
sp[4'd4][15][5] = 3'b111;\
sp[4'd4][15][6] = 3'b111;\
sp[4'd4][15][7] = 3'b111;\
sp[4'd4][15][8] = 3'b111;\
sp[4'd4][15][9] = 3'b111;\
sp[4'd4][15][10] = 3'b111;\
sp[4'd4][15][11] = 3'b111;\
sp[4'd4][15][12] = 3'b111;\
sp[4'd4][15][13] = 3'b111;\
sp[4'd4][15][14] = 3'b111;\
sp[4'd4][15][15] = 3'b111;

`define SNAKE_TAIL_PIC \
sp[4'd1][0][0] = 3'b111;\
sp[4'd1][0][1] = 3'b111;\
sp[4'd1][0][2] = 3'b111;\
sp[4'd1][0][3] = 3'b111;\
sp[4'd1][0][4] = 3'b111;\
sp[4'd1][0][5] = 3'b111;\
sp[4'd1][0][6] = 3'b111;\
sp[4'd1][0][7] = 3'b111;\
sp[4'd1][0][8] = 3'b111;\
sp[4'd1][0][9] = 3'b111;\
sp[4'd1][0][10] = 3'b111;\
sp[4'd1][0][11] = 3'b111;\
sp[4'd1][0][12] = 3'b111;\
sp[4'd1][0][13] = 3'b111;\
sp[4'd1][0][14] = 3'b111;\
sp[4'd1][0][15] = 3'b111;\
sp[4'd1][1][0] = 3'b111;\
sp[4'd1][1][1] = 3'b111;\
sp[4'd1][1][2] = 3'b111;\
sp[4'd1][1][3] = 3'b111;\
sp[4'd1][1][4] = 3'b111;\
sp[4'd1][1][5] = 3'b111;\
sp[4'd1][1][6] = 3'b111;\
sp[4'd1][1][7] = 3'b111;\
sp[4'd1][1][8] = 3'b111;\
sp[4'd1][1][9] = 3'b111;\
sp[4'd1][1][10] = 3'b111;\
sp[4'd1][1][11] = 3'b111;\
sp[4'd1][1][12] = 3'b111;\
sp[4'd1][1][13] = 3'b111;\
sp[4'd1][1][14] = 3'b111;\
sp[4'd1][1][15] = 3'b111;\
sp[4'd1][2][0] = 3'b111;\
sp[4'd1][2][1] = 3'b111;\
sp[4'd1][2][2] = 3'b111;\
sp[4'd1][2][3] = 3'b111;\
sp[4'd1][2][4] = 3'b111;\
sp[4'd1][2][5] = 3'b111;\
sp[4'd1][2][6] = 3'b111;\
sp[4'd1][2][7] = 3'b111;\
sp[4'd1][2][8] = 3'b111;\
sp[4'd1][2][9] = 3'b111;\
sp[4'd1][2][10] = 3'b111;\
sp[4'd1][2][11] = 3'b111;\
sp[4'd1][2][12] = 3'b111;\
sp[4'd1][2][13] = 3'b111;\
sp[4'd1][2][14] = 3'b111;\
sp[4'd1][2][15] = 3'b111;\
sp[4'd1][3][0] = 3'b111;\
sp[4'd1][3][1] = 3'b111;\
sp[4'd1][3][2] = 3'b111;\
sp[4'd1][3][3] = 3'b111;\
sp[4'd1][3][4] = 3'b000;\
sp[4'd1][3][5] = 3'b000;\
sp[4'd1][3][6] = 3'b000;\
sp[4'd1][3][7] = 3'b000;\
sp[4'd1][3][8] = 3'b000;\
sp[4'd1][3][9] = 3'b000;\
sp[4'd1][3][10] = 3'b000;\
sp[4'd1][3][11] = 3'b000;\
sp[4'd1][3][12] = 3'b111;\
sp[4'd1][3][13] = 3'b111;\
sp[4'd1][3][14] = 3'b111;\
sp[4'd1][3][15] = 3'b111;\
sp[4'd1][4][0] = 3'b111;\
sp[4'd1][4][1] = 3'b111;\
sp[4'd1][4][2] = 3'b111;\
sp[4'd1][4][3] = 3'b000;\
sp[4'd1][4][4] = 3'b000;\
sp[4'd1][4][5] = 3'b010;\
sp[4'd1][4][6] = 3'b010;\
sp[4'd1][4][7] = 3'b010;\
sp[4'd1][4][8] = 3'b010;\
sp[4'd1][4][9] = 3'b010;\
sp[4'd1][4][10] = 3'b010;\
sp[4'd1][4][11] = 3'b000;\
sp[4'd1][4][12] = 3'b000;\
sp[4'd1][4][13] = 3'b111;\
sp[4'd1][4][14] = 3'b111;\
sp[4'd1][4][15] = 3'b111;\
sp[4'd1][5][0] = 3'b111;\
sp[4'd1][5][1] = 3'b111;\
sp[4'd1][5][2] = 3'b111;\
sp[4'd1][5][3] = 3'b000;\
sp[4'd1][5][4] = 3'b010;\
sp[4'd1][5][5] = 3'b110;\
sp[4'd1][5][6] = 3'b110;\
sp[4'd1][5][7] = 3'b010;\
sp[4'd1][5][8] = 3'b010;\
sp[4'd1][5][9] = 3'b110;\
sp[4'd1][5][10] = 3'b110;\
sp[4'd1][5][11] = 3'b010;\
sp[4'd1][5][12] = 3'b000;\
sp[4'd1][5][13] = 3'b111;\
sp[4'd1][5][14] = 3'b111;\
sp[4'd1][5][15] = 3'b111;\
sp[4'd1][6][0] = 3'b111;\
sp[4'd1][6][1] = 3'b111;\
sp[4'd1][6][2] = 3'b111;\
sp[4'd1][6][3] = 3'b000;\
sp[4'd1][6][4] = 3'b010;\
sp[4'd1][6][5] = 3'b110;\
sp[4'd1][6][6] = 3'b001;\
sp[4'd1][6][7] = 3'b010;\
sp[4'd1][6][8] = 3'b010;\
sp[4'd1][6][9] = 3'b001;\
sp[4'd1][6][10] = 3'b110;\
sp[4'd1][6][11] = 3'b010;\
sp[4'd1][6][12] = 3'b000;\
sp[4'd1][6][13] = 3'b111;\
sp[4'd1][6][14] = 3'b111;\
sp[4'd1][6][15] = 3'b111;\
sp[4'd1][7][0] = 3'b111;\
sp[4'd1][7][1] = 3'b111;\
sp[4'd1][7][2] = 3'b111;\
sp[4'd1][7][3] = 3'b000;\
sp[4'd1][7][4] = 3'b010;\
sp[4'd1][7][5] = 3'b010;\
sp[4'd1][7][6] = 3'b010;\
sp[4'd1][7][7] = 3'b100;\
sp[4'd1][7][8] = 3'b100;\
sp[4'd1][7][9] = 3'b010;\
sp[4'd1][7][10] = 3'b010;\
sp[4'd1][7][11] = 3'b010;\
sp[4'd1][7][12] = 3'b000;\
sp[4'd1][7][13] = 3'b111;\
sp[4'd1][7][14] = 3'b111;\
sp[4'd1][7][15] = 3'b111;\
sp[4'd1][8][0] = 3'b111;\
sp[4'd1][8][1] = 3'b111;\
sp[4'd1][8][2] = 3'b111;\
sp[4'd1][8][3] = 3'b000;\
sp[4'd1][8][4] = 3'b010;\
sp[4'd1][8][5] = 3'b010;\
sp[4'd1][8][6] = 3'b010;\
sp[4'd1][8][7] = 3'b100;\
sp[4'd1][8][8] = 3'b100;\
sp[4'd1][8][9] = 3'b010;\
sp[4'd1][8][10] = 3'b010;\
sp[4'd1][8][11] = 3'b010;\
sp[4'd1][8][12] = 3'b000;\
sp[4'd1][8][13] = 3'b111;\
sp[4'd1][8][14] = 3'b111;\
sp[4'd1][8][15] = 3'b111;\
sp[4'd1][9][0] = 3'b111;\
sp[4'd1][9][1] = 3'b111;\
sp[4'd1][9][2] = 3'b111;\
sp[4'd1][9][3] = 3'b000;\
sp[4'd1][9][4] = 3'b010;\
sp[4'd1][9][5] = 3'b110;\
sp[4'd1][9][6] = 3'b001;\
sp[4'd1][9][7] = 3'b010;\
sp[4'd1][9][8] = 3'b010;\
sp[4'd1][9][9] = 3'b001;\
sp[4'd1][9][10] = 3'b110;\
sp[4'd1][9][11] = 3'b010;\
sp[4'd1][9][12] = 3'b000;\
sp[4'd1][9][13] = 3'b111;\
sp[4'd1][9][14] = 3'b111;\
sp[4'd1][9][15] = 3'b111;\
sp[4'd1][10][0] = 3'b111;\
sp[4'd1][10][1] = 3'b111;\
sp[4'd1][10][2] = 3'b111;\
sp[4'd1][10][3] = 3'b000;\
sp[4'd1][10][4] = 3'b010;\
sp[4'd1][10][5] = 3'b110;\
sp[4'd1][10][6] = 3'b110;\
sp[4'd1][10][7] = 3'b010;\
sp[4'd1][10][8] = 3'b010;\
sp[4'd1][10][9] = 3'b110;\
sp[4'd1][10][10] = 3'b110;\
sp[4'd1][10][11] = 3'b010;\
sp[4'd1][10][12] = 3'b000;\
sp[4'd1][10][13] = 3'b111;\
sp[4'd1][10][14] = 3'b111;\
sp[4'd1][10][15] = 3'b111;\
sp[4'd1][11][0] = 3'b111;\
sp[4'd1][11][1] = 3'b111;\
sp[4'd1][11][2] = 3'b111;\
sp[4'd1][11][3] = 3'b000;\
sp[4'd1][11][4] = 3'b000;\
sp[4'd1][11][5] = 3'b010;\
sp[4'd1][11][6] = 3'b010;\
sp[4'd1][11][7] = 3'b010;\
sp[4'd1][11][8] = 3'b010;\
sp[4'd1][11][9] = 3'b010;\
sp[4'd1][11][10] = 3'b010;\
sp[4'd1][11][11] = 3'b000;\
sp[4'd1][11][12] = 3'b000;\
sp[4'd1][11][13] = 3'b111;\
sp[4'd1][11][14] = 3'b111;\
sp[4'd1][11][15] = 3'b111;\
sp[4'd1][12][0] = 3'b111;\
sp[4'd1][12][1] = 3'b111;\
sp[4'd1][12][2] = 3'b111;\
sp[4'd1][12][3] = 3'b111;\
sp[4'd1][12][4] = 3'b000;\
sp[4'd1][12][5] = 3'b000;\
sp[4'd1][12][6] = 3'b000;\
sp[4'd1][12][7] = 3'b000;\
sp[4'd1][12][8] = 3'b000;\
sp[4'd1][12][9] = 3'b000;\
sp[4'd1][12][10] = 3'b000;\
sp[4'd1][12][11] = 3'b000;\
sp[4'd1][12][12] = 3'b111;\
sp[4'd1][12][13] = 3'b111;\
sp[4'd1][12][14] = 3'b111;\
sp[4'd1][12][15] = 3'b111;\
sp[4'd1][13][0] = 3'b111;\
sp[4'd1][13][1] = 3'b111;\
sp[4'd1][13][2] = 3'b111;\
sp[4'd1][13][3] = 3'b111;\
sp[4'd1][13][4] = 3'b111;\
sp[4'd1][13][5] = 3'b111;\
sp[4'd1][13][6] = 3'b111;\
sp[4'd1][13][7] = 3'b111;\
sp[4'd1][13][8] = 3'b111;\
sp[4'd1][13][9] = 3'b111;\
sp[4'd1][13][10] = 3'b111;\
sp[4'd1][13][11] = 3'b111;\
sp[4'd1][13][12] = 3'b111;\
sp[4'd1][13][13] = 3'b111;\
sp[4'd1][13][14] = 3'b111;\
sp[4'd1][13][15] = 3'b111;\
sp[4'd1][14][0] = 3'b111;\
sp[4'd1][14][1] = 3'b111;\
sp[4'd1][14][2] = 3'b111;\
sp[4'd1][14][3] = 3'b111;\
sp[4'd1][14][4] = 3'b111;\
sp[4'd1][14][5] = 3'b111;\
sp[4'd1][14][6] = 3'b111;\
sp[4'd1][14][7] = 3'b111;\
sp[4'd1][14][8] = 3'b111;\
sp[4'd1][14][9] = 3'b111;\
sp[4'd1][14][10] = 3'b111;\
sp[4'd1][14][11] = 3'b111;\
sp[4'd1][14][12] = 3'b111;\
sp[4'd1][14][13] = 3'b111;\
sp[4'd1][14][14] = 3'b111;\
sp[4'd1][14][15] = 3'b111;\
sp[4'd1][15][0] = 3'b111;\
sp[4'd1][15][1] = 3'b111;\
sp[4'd1][15][2] = 3'b111;\
sp[4'd1][15][3] = 3'b111;\
sp[4'd1][15][4] = 3'b111;\
sp[4'd1][15][5] = 3'b111;\
sp[4'd1][15][6] = 3'b111;\
sp[4'd1][15][7] = 3'b111;\
sp[4'd1][15][8] = 3'b111;\
sp[4'd1][15][9] = 3'b111;\
sp[4'd1][15][10] = 3'b111;\
sp[4'd1][15][11] = 3'b111;\
sp[4'd1][15][12] = 3'b111;\
sp[4'd1][15][13] = 3'b111;\
sp[4'd1][15][14] = 3'b111;\
sp[4'd1][15][15] = 3'b111;

`define SPRITE_INIT `APPLE_PIC `SNAKE_HEAD_PIC `SNAKE_TAIL_PIC

`endif // sprites_vh
