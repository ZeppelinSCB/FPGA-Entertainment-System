module letter_game_won
(
    letter_x        ,
    letter_y        ,
    letter_won    ,
    letter_won_o        
);

input   [7:0]   letter_x     ;//x coordinate of pixel with respect to letter
input   [7:0]   letter_y     ;//y coordinate of pixel with respect to letter

output  [0:0]   letter_won_o     ;//letter output


assign          letter_won[ 0] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[ 1] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[ 2] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[ 3] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[ 4] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[ 5] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[ 6] <= {8'b00000000, 8'b11111110, 8'b00111111, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b11111110, 8'b01111111, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111110, 8'b01111111, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b11111110, 8'b00111111, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11100000, 8'b00000000};
assign          letter_won[ 7] <= {8'b00000000, 8'b01111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b01111011, 8'b11011110, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b11111100, 8'b00000000, 8'b00000000, 8'b01111100, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b01111100, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01111110, 8'b00000000, 8'b00000000, 8'b01111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01111110, 8'b00000000, 8'b00000000, 8'b01111101, 8'b11111000, 8'b00000000};
assign          letter_won[ 8] <= {8'b00000000, 8'b00111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00011110, 8'b00000000, 8'b00000000, 8'b01110011, 8'b11001110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00011110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b01111100, 8'b00000000};
assign          letter_won[ 9] <= {8'b00000000, 8'b00111100, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b11100011, 8'b11000110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00111100, 8'b00000000};
assign          letter_won[10] <= {8'b00000000, 8'b00111100, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b11100011, 8'b11000111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00011100, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_won[11] <= {8'b00000000, 8'b00111100, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_won[12] <= {8'b00000000, 8'b00011100, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00011110, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001110, 8'b11100000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00011100, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_won[13] <= {8'b00000000, 8'b00011110, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00001111, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001110, 8'b11100000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00111000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001110, 8'b00000000};
assign          letter_won[14] <= {8'b00000000, 8'b00011110, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00001111, 8'b01100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001110, 8'b11110000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_won[15] <= {8'b00000000, 8'b00011110, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00111100, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00001100, 8'b11110000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00011110, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_won[16] <= {8'b00000000, 8'b00001110, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011100, 8'b01110000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00001110, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_won[17] <= {8'b00000000, 8'b00001110, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00111101, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011100, 8'b01110000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00001110, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_won[18] <= {8'b00000000, 8'b00001111, 8'b01100000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00111101, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011100, 8'b01111000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b01100000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_won[19] <= {8'b00000000, 8'b00001111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00111100, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00001111, 8'b00000000};
assign          letter_won[20] <= {8'b00000000, 8'b00001111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00001111, 8'b00000000, 8'b00000000, 8'b00111100, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b01111000, 8'b00000000, 8'b00000000, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11100000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00110000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_won[21] <= {8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01110000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00111000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_won[22] <= {8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000111, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000011, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000011, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_won[23] <= {8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011110, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01111000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00110000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00000110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000111, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00011110, 8'b00000000};
assign          letter_won[24] <= {8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00000111, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00000110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b00111100, 8'b00000000};
assign          letter_won[25] <= {8'b00000000, 8'b00000011, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111110, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b01110000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00111110, 8'b00011100, 8'b00000000, 8'b00000000, 8'b01111000, 8'b00011100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00001110, 8'b00000000, 8'b00000000, 8'b00111000, 8'b01111000, 8'b00000000};
assign          letter_won[26] <= {8'b00000000, 8'b00000011, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b11111000, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00011111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b01111100, 8'b00111110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b11000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01111110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00111100, 8'b01111110, 8'b00000000, 8'b00000000, 8'b01111111, 8'b11111000, 8'b00000000};
assign          letter_won[27] <= {8'b00000000, 8'b00000011, 8'b10000000, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b00011111, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000001, 8'b11111100, 8'b01111111, 8'b00000000, 8'b00000000, 8'b00001111, 8'b11110000, 8'b00000000, 8'b00000000, 8'b11111110, 8'b01111111, 8'b00000000, 8'b00000000, 8'b00111111, 8'b11111100, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b00000011, 8'b10000000, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11111110, 8'b00000000, 8'b00000000, 8'b11111111, 8'b11100000, 8'b00000000};
assign          letter_won[28] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[29] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[30] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
assign          letter_won[31] <= {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};


always@(*)
begin
    letter_won_o = letter_won[letter_y][letter_x];
end

endmodule