`include "../libs/define.vh"

module key_in
(
    key_up          , 
    key_down        , 
    key_left        , 
    key_right       ,
    key_flag        , 
    iClk             ,
    sys_clk         ,
    sys_rst_n       ,
    oDirection

);

input wire key_up        ;//key1
input wire key_down      ;//key2
input wire key_left      ;//key0
input wire key_right     ;//key3
input wire key_flag		 ;
input wire iClk          ;
input wire sys_clk       ;
input wire sys_rst_n     ;

output reg [0:1] oDirection;


reg left, right, up, down;
reg key_press;
reg [19:0] cnt_20ms ;

parameter CNT_MAX = 20'd999_999;//The maximum counter number

initial

begin
    oDirection = `TOP_DIR;
end

always @(posedge sys_clk or negedge sys_rst_n) begin

    key_press = (key_up||key_down||key_left||key_right);

 	if(sys_rst_n == 1'b0)
		cnt_20ms <= 20'b0;
	else if(key_press == 1'b1)
		cnt_20ms <= 20'b0;
	else if(cnt_20ms == CNT_MAX && key_press == 1'b0)
		cnt_20ms <= cnt_20ms;
	else
		cnt_20ms <= cnt_20ms + 1'b1;
end

always@(posedge sys_clk or negedge sys_rst_n) begin
	if(sys_rst_n == 1'b0)
		key_flag <= 1'b0;
	else if(cnt_20ms == CNT_MAX - 1'b1)
		key_flag <= 1'b1;
	else
		key_flag <= 1'b0;
end

always @(posedge iClk)
begin

    left = key_left		;//left = two_resistors_x;
    right = key_right	;//right = ~one_resistor_x;
    up = key_up			;//up = two_resistors_y;
    down = key_down		;//down = ~one_resistor_y;

	if((left + right + up + down == 3'b001)&&(key_flag == 1'b1)) // if only one pressed 

	begin 

		if(left && (oDirection != `RIGHT_DIR)) 

		begin 
			oDirection = `LEFT_DIR; 
		end 



		if(right && (oDirection != `LEFT_DIR)) 

		begin 
			oDirection = `RIGHT_DIR; 
		end 



		if(up && (oDirection != `DOWN_DIR)) 

		begin 
			oDirection = `TOP_DIR;
		end 			 



		if(down && (oDirection != `TOP_DIR)) 

		begin 
			oDirection = `DOWN_DIR; 
		end 
	end

    else
        oDirection = oDirection; 

end

endmodule