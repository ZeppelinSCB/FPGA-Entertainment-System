/*

*/
Map_Hori
Map_Vert

module Tile_Renderer(
    input wire sys_clk,
    input wire sys_rst_n,
    input wire tile_map_rom,
    
)

endmodule